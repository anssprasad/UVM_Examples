//------------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//   
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//   
//       http://www.apache.org/licenses/LICENSE-2.0
//   
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

//----------------------------------------------------------------------
//   THIS IS AUTOMATICALLY GENERATED CODE
//   Generated by Mentor Graphics' Register Assistant V2010.1 (Build 2) Beta
//   UVM Register Kit version 2.0
//----------------------------------------------------------------------
// Project         : wb_registers
// Unit            : wb_register_pkg
// File            : wb_register_pkg.sv
//----------------------------------------------------------------------
// Created by      : mike
// Creation Date   : 6/1/10 10:59 AM
//----------------------------------------------------------------------
// Title           : wb_registers
//
// Description     : 
//
//----------------------------------------------------------------------

//----------------------------------------------------------------------
// wb_register_pkg
//----------------------------------------------------------------------
package wb_register_pkg;

  import uvm_pkg::*;
  import uvm_register_pkg::*;
  `include "uvm_register_macros.svh" // -*- FIXME include of uvm file other than uvm_macros.svh detected, you should move to an import based methodology
  
  /* DEFINE TYPES FOR THE DATA CONTAINED IN THE REGISTERS */
  
  // Types for enums


  // Types for non-field registers

   typedef bit[31:0] bit32_t;


  // Types for registers which have fields


   typedef struct packed {
      // reserved bit field
      bit[31:17] reserved;
      // Receive Small
      bit rec_small;
      // Pad Enable 
      bit pad;
      // Huge Enable 
      bit huge_en;
      // CRC Enable 
      bit crc_en;
      // Delayed CRC Enable 
      bit dly_crc_en;
      // Reset MAC 
      bit rst;
      // Full Duplex 
      bit full_d;
      // Excess Defer 
      bit ex_defer;
      // No Backoff 
      bit no_back_off;
      // Loop Back 
      bit loop_back;
      // Min. IFG not required 
      bit ifg;
      // Promiscuous (receive all)
      bit pro;
      // Use Individual Hash 
      bit iam;
      // Reject Broadcast
      bit bro;
      // No Preamble 
      bit nopre;
      // Transmit Enable 
      bit txen;
      // Receive Enable  
      bit rxen;
   } mode_register_t;

   typedef struct packed {
      // reserved bit field
      bit[31:7] reserved;
      // Receive control frame 
      bit rxc;
      // Transmit Control Frame
      bit txc;
      // Busy mask 
      bit busy;
      // Receive error 
      bit rxe;
      // receive frame 
      bit rxb;
      // transmit error 
      bit txe;
      // Transmit buffer   
      bit txb;
   } irq_source_register_t;

   typedef struct packed {
      // reserved bit field   
      bit[31:7] reserved;
      // Receive control frame mask 
      bit rxc_m;
      // Transmit Control Frame mask
      bit txc_m;
      // Busy mask 
      bit busy_m;
      // Receive error mask
      bit rxe_m;
      // receive frame mask
      bit rxb_m;
      // transmit error mask
      bit txe_m;
      // Transmit buffer mask  
      bit txb_m;
   } int_mask_register_t;

   typedef struct packed {
      // Tx BD length 
      bit[31:16] len;
      // Tx BD Ready 
      bit rdy;
      // Tx BD IRQ Enable
      bit irq;
      // Tx BD Wrap (last BD) 
      bit wrap;
      // Tx BD Pad Enable 
      bit pad_en;
      // Tx BD CRC Enable
      bit crc_en;
      // reserved bit field
      bit[10:9] reserved;
      // Tx BD Underrun Status 
      bit under_run;
      // Tx BD Retry Status 
      bit[7:4] retry;
      // Tx BD Retransmission Limit Status 
      bit ret_lim;
      // Tx BD Late Collision Status 
      bit late_col;
      // Tx BD Defer Status 
      bit defer;
      // Tx BD Carrier Sense Lost Status 
      bit c_sense;
   } tx_bd_t;

   typedef struct packed {
      // Rx BD length 
      bit[31:16] len;
      // Rx BD Ready 
      bit rdy;
      // Rx BD IRQ Enable
      bit irq;
      // Rx BD Wrap (last BD) 
      bit wrap;
      // reserved bit field
      bit[12:9] reserved;
      // Rx BD Control frame 
      bit c_frame;
      // Rx BD Miss Status 
      bit miss;
      // Rx BD Overrun Status 
      bit over_run;
      // Rx BD Invalid Symbol Status 
      bit inval_symbol;
      // Rx BD Dribble Nibble Status 
      bit dn;
      // Rx BD Too Long Status 
      bit too_long;
      // Rx BD Too Short Frame Status
      bit s_frame;
      // Rx BD CRC Error Status 
      bit crc_error;
      // Rx BD Late Collision Status 
      bit l_coll;
   } rx_bd_t;




  /* DEFINE REGISTER CLASSES */



   //--------------------------------------------------------------------
   // rx_bd_ptr
   //--------------------------------------------------------------------
   // RX BD Pointer
   class rx_bd_ptr extends uvm_register #(bit32_t);
      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         
      endfunction
   endclass
   //--------------------------------------------------------------------
   // mac_addr0_register
   //--------------------------------------------------------------------
   // MAC Addr0 Register
   class mac_addr0_register extends uvm_register #(bit32_t);
      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         
      endfunction
   endclass

   //--------------------------------------------------------------------
   // irq_source_register
   //--------------------------------------------------------------------
   // IRQ Source Register
   class irq_source_register extends uvm_register #(irq_source_register_t);
      `uvm_register_begin_fields
         `uvm_register_field(rxc)
         `uvm_register_field(txc)
         `uvm_register_field(busy)
         `uvm_register_field(rxe)
         `uvm_register_field(rxb)
         `uvm_register_field(txe)
         `uvm_register_field(txb)
      `uvm_register_end_fields

      //--------------------------------------------------------------------
      // coverage
      //--------------------------------------------------------------------
      covergroup c;
         rxc    : coverpoint data.rxc;
         txc    : coverpoint data.txc;
         busy   : coverpoint data.busy;
         rxe    : coverpoint data.rxe;
         rxb    : coverpoint data.rxb;
         txe    : coverpoint data.txe;
         txb    : coverpoint data.txb;
      endgroup
      //--------------------------------------------------------------------
      // sample
      //--------------------------------------------------------------------
      function void sample();
         c.sample();
      endfunction

      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         c = new();

         uvm_report_info("irq_source_register", "new()");
         add_field("rxc",  1'b0, "W1C");
         add_field("txc",  1'b0, "W1C");
         add_field("busy", 1'b0, "W1C");
         add_field("rxe",  1'b0, "W1C");
         add_field("rxb",  1'b0, "W1C");
         add_field("txe",  1'b0, "W1C");
         add_field("txb",  1'b0, "W1C");
      endfunction

      //--------------------------------------------------------------------
      // convert2string
      //--------------------------------------------------------------------
      function string convert2string();
         return $psprintf("CSR: (%p) (%x %x %x %x %x %x %x %x )", data, data.reserved, data.rxc, data.txc, data.busy, data.rxe, data.rxb, data.txe, data.txb);
      endfunction
   endclass


   //--------------------------------------------------------------------
   // mode_register
   //--------------------------------------------------------------------
   // Mode Register
   class mode_register extends uvm_register #(mode_register_t);
      `uvm_register_begin_fields
         `uvm_register_field(rec_small)
         `uvm_register_field(pad)
         `uvm_register_field(huge_en)
         `uvm_register_field(crc_en)
         `uvm_register_field(dly_crc_en)
         `uvm_register_field(rst)
         `uvm_register_field(full_d)
         `uvm_register_field(ex_defer)
         `uvm_register_field(no_back_off)
         `uvm_register_field(loop_back)
         `uvm_register_field(ifg)
         `uvm_register_field(pro)
         `uvm_register_field(iam)
         `uvm_register_field(bro)
         `uvm_register_field(nopre)
         `uvm_register_field(txen)
         `uvm_register_field(rxen)
      `uvm_register_end_fields

      //--------------------------------------------------------------------
      // coverage
      //--------------------------------------------------------------------
      covergroup c;
         rec_small    : coverpoint data.rec_small;
         pad    : coverpoint data.pad;
         huge_en   : coverpoint data.huge_en;
         crc_en    : coverpoint data.crc_en;
         dly_crc_en   : coverpoint data.dly_crc_en;
         rst    : coverpoint data.rst;
         full_d    : coverpoint data.full_d;
         ex_defer  : coverpoint data.ex_defer;
         no_back_off  : coverpoint data.no_back_off;
         loop_back    : coverpoint data.loop_back;
         ifg    : coverpoint data.ifg;
         pro    : coverpoint data.pro;
         iam    : coverpoint data.iam;
         bro    : coverpoint data.bro;
         nopre  : coverpoint data.nopre;
         txen   : coverpoint data.txen;
         rxen   : coverpoint data.rxen;
      endgroup
      //--------------------------------------------------------------------
      // sample
      //--------------------------------------------------------------------
      function void sample();
         c.sample();
      endfunction

      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         c = new();

         uvm_report_info("mode_register", "new()");
         add_field("rec_small",  1'b0, "RW");
         add_field("pad",  1'b1, "RW");
         add_field("huge_en", 1'b0, "RW");
         add_field("crc_en",  1'b1, "RW");
         add_field("dly_crc_en", 1'b0, "RW");
         add_field("rst",  1'b0, "RW");
         add_field("full_d",  1'b0, "RW");
         add_field("ex_defer",   1'b0, "RW");
         add_field("no_back_off",   1'b0, "RW");
         add_field("loop_back",  1'b0, "RW");
         add_field("ifg",  1'b0, "RW");
         add_field("pro",  1'b0, "RW");
         add_field("iam",  1'b0, "RW");
         add_field("bro",  1'b0, "RW");
         add_field("nopre",   1'b0, "RW");
         add_field("txen", 1'b1, "RW");
         add_field("rxen", 1'b0, "RW");
      endfunction

      //--------------------------------------------------------------------
      // convert2string
      //--------------------------------------------------------------------
      function string convert2string();
         return $psprintf("CSR: (%p) (%x %x %x %x %x %x %x %x %x %x %x %x %x %x %x %x %x %x )", data, data.reserved, data.rec_small, data.pad, data.huge_en, data.crc_en, data.dly_crc_en, data.rst, data.full_d, data.ex_defer, data.no_back_off, data.loop_back, data.ifg, data.pro, data.iam, data.bro, data.nopre, data.txen, data.rxen);
      endfunction
   endclass

   //--------------------------------------------------------------------
   // mac_addr1_register
   //--------------------------------------------------------------------
   // MAC Addr1 Register
   class mac_addr1_register extends uvm_register #(bit32_t);
      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         
      endfunction
   endclass

   //--------------------------------------------------------------------
   // rx_bd
   //--------------------------------------------------------------------
   // RX Buffer Descriptor
   class rx_bd extends uvm_register #(rx_bd_t);
      `uvm_register_begin_fields
         `uvm_register_field(len)
         `uvm_register_field(rdy)
         `uvm_register_field(irq)
         `uvm_register_field(wrap)
         `uvm_register_field(c_frame)
         `uvm_register_field(miss)
         `uvm_register_field(over_run)
         `uvm_register_field(inval_symbol)
         `uvm_register_field(dn)
         `uvm_register_field(too_long)
         `uvm_register_field(s_frame)
         `uvm_register_field(crc_error)
         `uvm_register_field(l_coll)
      `uvm_register_end_fields

      //--------------------------------------------------------------------
      // coverage
      //--------------------------------------------------------------------
      covergroup c;
         len    : coverpoint data.len;
         rdy    : coverpoint data.rdy;
         irq    : coverpoint data.irq;
         wrap   : coverpoint data.wrap;
         c_frame   : coverpoint data.c_frame;
         miss   : coverpoint data.miss;
         over_run  : coverpoint data.over_run;
         inval_symbol    : coverpoint data.inval_symbol;
         dn  : coverpoint data.dn;
         too_long  : coverpoint data.too_long;
         s_frame   : coverpoint data.s_frame;
         crc_error    : coverpoint data.crc_error;
         l_coll    : coverpoint data.l_coll;
      endgroup
      //--------------------------------------------------------------------
      // sample
      //--------------------------------------------------------------------
      function void sample();
         c.sample();
      endfunction

      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         c = new();

         uvm_report_info("rx_bd", "new()");
         add_field("len",  16'h0000,   "RW");
         add_field("rdy",  1'b1, "RW");
         add_field("irq",  1'b0, "RW");
         add_field("wrap", 1'b1, "RW");
         add_field("c_frame", 1'b1, "RW");
         add_field("miss", 1'b0, "RW");
         add_field("over_run",   1'b1, "RW");
         add_field("inval_symbol",  1'b0, "RW");
         add_field("dn",   1'b1, "RW");
         add_field("too_long",   1'b0, "RW");
         add_field("s_frame", 1'b1, "RW");
         add_field("crc_error",  1'b0, "RW");
         add_field("l_coll",  1'b1, "RW");
      endfunction

      //--------------------------------------------------------------------
      // convert2string
      //--------------------------------------------------------------------
      function string convert2string();
         return $psprintf("CSR: (%p) (%x %x %x %x %x %x %x %x %x %x %x %x %x %x )", data, data.len, data.rdy, data.irq, data.wrap, data.reserved, data.c_frame, data.miss, data.over_run, data.inval_symbol, data.dn, data.too_long, data.s_frame, data.crc_error, data.l_coll);
      endfunction
   endclass


   //--------------------------------------------------------------------
   // int_mask_register
   //--------------------------------------------------------------------
   // IRQ Mask Register
   class int_mask_register extends uvm_register #(int_mask_register_t);
      `uvm_register_begin_fields
         `uvm_register_field(rxc_m)
         `uvm_register_field(txc_m)
         `uvm_register_field(busy_m)
         `uvm_register_field(rxe_m)
         `uvm_register_field(rxb_m)
         `uvm_register_field(txe_m)
         `uvm_register_field(txb_m)
      `uvm_register_end_fields

      //--------------------------------------------------------------------
      // coverage
      //--------------------------------------------------------------------
      covergroup c;
         rxc_m  : coverpoint data.rxc_m;
         txc_m  : coverpoint data.txc_m;
         busy_m    : coverpoint data.busy_m;
         rxe_m  : coverpoint data.rxe_m;
         rxb_m  : coverpoint data.rxb_m;
         txe_m  : coverpoint data.txe_m;
         txb_m  : coverpoint data.txb_m;
      endgroup
      //--------------------------------------------------------------------
      // sample
      //--------------------------------------------------------------------
      function void sample();
         c.sample();
      endfunction

      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         c = new();

         uvm_report_info("int_mask_register", "new()");
         add_field("rxc_m",   1'b0, "RW");
         add_field("txc_m",   1'b0, "RW");
         add_field("busy_m",  1'b0, "RW");
         add_field("rxe_m",   1'b0, "RW");
         add_field("rxb_m",   1'b0, "RW");
         add_field("txe_m",   1'b0, "RW");
         add_field("txb_m",   1'b0, "RW");
      endfunction

      //--------------------------------------------------------------------
      // convert2string
      //--------------------------------------------------------------------
      function string convert2string();
         return $psprintf("CSR: (%p) (%x %x %x %x %x %x %x %x )", data, data.reserved, data.rxc_m, data.txc_m, data.busy_m, data.rxe_m, data.rxb_m, data.txe_m, data.txb_m);
      endfunction
   endclass


   //--------------------------------------------------------------------
   // tx_bd
   //--------------------------------------------------------------------
   // TX Buffer Descriptor
   class tx_bd extends uvm_register #(tx_bd_t);
      `uvm_register_begin_fields
         `uvm_register_field(len)
         `uvm_register_field(rdy)
         `uvm_register_field(irq)
         `uvm_register_field(wrap)
         `uvm_register_field(pad_en)
         `uvm_register_field(crc_en)
         `uvm_register_field(under_run)
         `uvm_register_field(retry)
         `uvm_register_field(ret_lim)
         `uvm_register_field(late_col)
         `uvm_register_field(defer)
         `uvm_register_field(c_sense)
      `uvm_register_end_fields

      //--------------------------------------------------------------------
      // coverage
      //--------------------------------------------------------------------
      covergroup c;
         len    : coverpoint data.len;
         rdy    : coverpoint data.rdy;
         irq    : coverpoint data.irq;
         wrap   : coverpoint data.wrap;
         pad_en    : coverpoint data.pad_en;
         crc_en    : coverpoint data.crc_en;
         under_run    : coverpoint data.under_run;
         retry  : coverpoint data.retry;
         ret_lim   : coverpoint data.ret_lim;
         late_col  : coverpoint data.late_col;
         defer  : coverpoint data.defer;
         c_sense   : coverpoint data.c_sense;
      endgroup
      //--------------------------------------------------------------------
      // sample
      //--------------------------------------------------------------------
      function void sample();
         c.sample();
      endfunction

      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         c = new();

         uvm_report_info("tx_bd", "new()");
         add_field("len",  16'h0000,   "RW");
         add_field("rdy",  1'b0, "RW");
         add_field("irq",  1'b0, "RW");
         add_field("wrap", 1'b0, "RW");
         add_field("pad_en",  1'b0, "RW");
         add_field("crc_en",  1'b0, "RW");
         add_field("under_run",  1'b0, "RW");
         add_field("retry",   4'h0, "RW");
         add_field("ret_lim", 1'b0, "RW");
         add_field("late_col",   1'b0, "RW");
         add_field("defer",   1'b0, "RW");
         add_field("c_sense", 1'b0, "RW");
      endfunction

      //--------------------------------------------------------------------
      // convert2string
      //--------------------------------------------------------------------
      function string convert2string();
         return $psprintf("CSR: (%p) (%x %x %x %x %x %x %x %x %x %x %x %x %x )", data, data.len, data.rdy, data.irq, data.wrap, data.pad_en, data.crc_en, data.reserved, data.under_run, data.retry, data.ret_lim, data.late_col, data.defer, data.c_sense);
      endfunction
   endclass

   //--------------------------------------------------------------------
   // tx_bd_ptr
   //--------------------------------------------------------------------
   // TX BD pointer
   class tx_bd_ptr extends uvm_register #(bit32_t);
      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         
      endfunction
   endclass


  /* REGISTER FILE */
   //--------------------------------------------------------------------
   // mac_reg_file
   //--------------------------------------------------------------------
   class mac_reg_file extends uvm_register_file;
      // mode reg instance
      mode_register  mode_reg;
      // irq source instance
      irq_source_register  irq_source_reg;
      // Int mask instance
      int_mask_register int_mask_reg;
      // MAC Addr 0 instance
      mac_addr0_register   mac_addr0_reg;
      // MAC Addr1 instance
      mac_addr1_register   mac_addr1_reg;
      // TX Buffer Descriptor 0
      tx_bd tx_bd_0;
      // TX Buffer Descriptor 0 Ptr
      tx_bd_ptr   tx_bd_0_ptr;
      // RX Buffer Descriptor 0
      rx_bd rx_bd_0;
      // RX Buffer Descriptor 0 Ptr
      rx_bd_ptr   rx_bd_0_ptr;

      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
         uvm_report_info("mac_reg_file", "new()");

         mode_reg = new("mode_reg", this);
         irq_source_reg = new("irq_source_reg", this);
         int_mask_reg   = new("int_mask_reg", this);
         mac_addr0_reg  = new("mac_addr0_reg", this);
         mac_addr1_reg  = new("mac_addr1_reg", this);
         tx_bd_0  = new("tx_bd_0", this);
         tx_bd_0_ptr = new("tx_bd_0_ptr", this);
         rx_bd_0  = new("rx_bd_0", this);
         rx_bd_0_ptr = new("rx_bd_0_ptr", this);

         mode_reg.set_reset_value(32'h0000a002);
         irq_source_reg.set_reset_value(32'h00000000);
         int_mask_reg.set_reset_value(32'h00000000);
         mac_addr0_reg.set_reset_value(32'h00000000);
         mac_addr1_reg.set_reset_value(32'h00000000);
         tx_bd_0.set_reset_value(32'h00000000);
         tx_bd_0_ptr.set_reset_value(32'h00000000);
         rx_bd_0.set_reset_value(32'h00000001);
         rx_bd_0_ptr.set_reset_value(32'h00000002);

         add_register(mode_reg.get_fullname(),  'h00, mode_reg);
         add_register(irq_source_reg.get_fullname(),  'h04, irq_source_reg);
         add_register(int_mask_reg.get_fullname(), 'h08, int_mask_reg);
         add_register(mac_addr0_reg.get_fullname(),   'h40, mac_addr0_reg);
         add_register(mac_addr1_reg.get_fullname(),   'h44, mac_addr1_reg);
         add_register(tx_bd_0.get_fullname(),   'h400,   tx_bd_0);
         add_register(tx_bd_0_ptr.get_fullname(),  'h404,   tx_bd_0_ptr);
         add_register(rx_bd_0.get_fullname(),   'h600,   rx_bd_0);
         add_register(rx_bd_0_ptr.get_fullname(),  'h604,   rx_bd_0_ptr);

      endfunction
   endclass




  /* REGISTER MAP */
   //--------------------------------------------------------------------
   // wb_mem_map
   //--------------------------------------------------------------------
   class wb_mem_map extends uvm_register_map;
      // Registers for MAC 0
      mac_reg_file mac_0_regs;

      //--------------------------------------------------------------------
      // new
      //--------------------------------------------------------------------
      function new(string name, uvm_named_object parent);
         super.new(name, parent);
      endfunction
      //--------------------------------------------------------------------
      // build_maps
      //--------------------------------------------------------------------
      virtual function void build_maps();
         uvm_report_info("wb_mem_map", "build_maps()");

         //--------------------------------------------------------------------
         // Construct the instances
         //--------------------------------------------------------------------
         mac_0_regs = new("mac_0_regs", this);


         add_register_file(mac_0_regs, 32'h00100000);

      endfunction
   endclass

  //
  // Class to automatically load a register map.
  
  //----------------------------------------------------------------------
  // register_map_auto_load
  //----------------------------------------------------------------------
  class register_map_auto_load;

    // Triggers factory registration of this default
    //  sequence. Can be overriden by the user using
    //  "default_auto_register_test".
    register_sequence_all_registers
      #(uvm_register_transaction, 
        uvm_register_transaction) dummy;

    static bit loaded = build_register_map();

    static function bit build_register_map();

      wb_mem_map register_map;

      register_map = new("register_map", null);

      register_map.build_maps();

      uvm_config_db #(uvm_register_map)::set(null, "*","register_map", register_map);
      return 1;
    endfunction

  endclass
endpackage
