//
//------------------------------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------
//
// Package contains a simple env containing the mbus_agent
// and the mbus_test
//
package mbus_pipelined_env_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import mbus_pipelined_agent_pkg::*;

class mbus_pipelined_env extends uvm_component;

`uvm_component_utils(mbus_pipelined_env)

function new(string name = "mbus_pipelined_env", uvm_component parent = null);
  super.new(name, parent);
endfunction

mbus_pipelined_agent m_mbus_agent;

function void build_phase(uvm_phase phase);
  m_mbus_agent = mbus_pipelined_agent::type_id::create("m_bus_agent", this);
endfunction: build_phase

endclass: mbus_pipelined_env

class mbus_test extends uvm_test;

`uvm_component_utils(mbus_test)

function new(string name = "mbus_test", uvm_component parent = null);
  super.new(name, parent);
endfunction

// Need to be here since they contain check data
mbus_unpipelined_seq t_seq_1;
mbus_pipelined_seq t_seq_2;
mbus_pipelined_check_seq t_seq_3;
mbus_pipelined_check_rsp_handler_seq t_seq_4;


mbus_pipelined_env m_env;
mbus_pipelined_agent_config mbus_agent_cfg;

function void build_phase(uvm_phase phase);
  set_config_int("*", "recording_detail", UVM_FULL);
  mbus_agent_cfg =  mbus_pipelined_agent_config::type_id::create("mbus_agent_cfg");
  if (!uvm_config_db #(virtual mbus_if)::get(this, "", "MBUS_vif", mbus_agent_cfg.MBUS)) begin
    `uvm_error("Build", "MBUS_vif not found")
  end
  uvm_config_db #(mbus_pipelined_agent_config)::set(this, "*", "mbus_agent_config", mbus_agent_cfg);
  m_env = mbus_pipelined_env::type_id::create("menv", this);
endfunction: build_phase

task run_phase(uvm_phase phase);

  phase.raise_objection(this, "Starting test");
  t_seq_1 = mbus_unpipelined_seq::type_id::create("t_seq_1");
  t_seq_2 = mbus_pipelined_seq::type_id::create("t_seq_2");
  t_seq_3 = mbus_pipelined_check_seq::type_id::create("t_seq_3");
  t_seq_3.base_address = 32'h0010_0000;
  t_seq_4 = mbus_pipelined_check_rsp_handler_seq::type_id::create("t_seq_4");
  t_seq_4.base_address = 32'h0012_0000;


  t_seq_1.start(m_env.m_mbus_agent.m_sequencer);
  t_seq_2.start(m_env.m_mbus_agent.m_sequencer);
  fork
    t_seq_1.start(m_env.m_mbus_agent.m_sequencer);
    t_seq_2.start(m_env.m_mbus_agent.m_sequencer);
  join
  phase.drop_objection(this, "Ending test");
endtask: run_phase

function void report_phase(uvm_phase phase);
  if((t_seq_1.error_count == 0) && (t_seq_3.error_count == 0) && (t_seq_4.error_count == 0)) begin
    `uvm_info("** UVM TEST PASSED **", "No errors occurred", UVM_LOW)
  end
  else begin
    `uvm_error("** UVM TEST FAILED **", "Errors occurred")
  end
endfunction: report_phase

endclass: mbus_test
/*
class mbus_test_c extends uvm_test;

`uvm_component_utils(mbus_test_c)

function new(string name = "mbus_test_c", uvm_component parent = null);
  super.new(name, parent);
endfunction

mbus_pipelined_env m_env;
mbus_pipelined_agent_config mbus_agent_cfg;

function void build_phase(uvm_phase phase);
  set_config_int("*", "recording_detail", UVM_FULL);
  mbus_agent_cfg =  mbus_pipelined_agent_config::type_id::create("mbus_agent_cfg");
  if (!uvm_config_db #(virtual mbus_if)::get(this, "", "MBUS_vif", mbus_agent_cfg.MBUS)) begin
    `uvm_error("Build", "MBUS_vif not found")
  end
  uvm_config_db #(mbus_pipelined_agent_config)::set(this, "*", "mbus_agent_config", mbus_agent_cfg);
  m_env = mbus_pipelined_env::type_id::create("menv", this);
endfunction: build_phase

task run_phase(uvm_phase phase);
  mbus_complete_trans_seq t_seq_1;

  phase.raise_objection(this, "Starting test");
  t_seq_1 = mbus_complete_trans_seq::type_id::create("t_seq_1");
  t_seq_1.start_address = 32'h0012_0000;

  fork
    t_seq_1.start(m_env.m_mbus_agent.m_sequencer);
  join
  phase.drop_objection(this, "Ending test");
endtask: run_phase

endclass: mbus_test_c
*/
endpackage: mbus_pipelined_env_pkg

module top_tb;

import uvm_pkg::*;
import mbus_pipelined_env_pkg::*;

mbus_if MBUS();
gpio_if GPIO();

mbus_slave dut(.bus(MBUS), .gpio(GPIO));

// Clock and reset process
initial
  begin
    MBUS.MRESETN = 0;
    MBUS.MCLK = 0;
    repeat(6) begin
      #10 MBUS.MCLK = ~MBUS.MCLK;
    end
    MBUS.MRESETN = 1;
    forever begin
      #10 MBUS.MCLK = ~MBUS.MCLK;
    end
  end

// GPIO Clock
assign GPIO.clk = MBUS.MCLK;

// UVM Starting process
initial
  begin
    // Setup the virtual interfaces
    uvm_config_db #(virtual mbus_if)::set(null, "uvm_test_top", "MBUS_vif" , MBUS);
    uvm_config_db #(virtual gpio_if)::set(null, "uvm_test_top", "GPIO_vif" , GPIO);
    // Start up the uvm test bench
    run_test("mbus_test");
  end

endmodule: top_tb
