//------------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

module top_hdl;

`include "timescale.v"

// PCLK and PRESETn
//
logic PCLK;
logic PRESETn;

//
// Instantiate the interfaces:
//
apb_if APB(PCLK, PRESETn);  // APB interface
spi_if SPI(PCLK, PRESETN);  // SPI Interface

intr_if INTR(PCLK, PRESETn);   // Interrupt

// tbx vif_binding_block
initial begin
  import uvm_pkg::uvm_config_db;
  uvm_config_db #(virtual intr_if) C;
  C.set(null, "uvm_test_top", $psprintf("%m.INTR") , INTR);
end

//if(HAS_APB_AGENT) begin: has_apb_agent
apb_driver_bfm  APB_DRIVER(APB.driver_mp);
apb_monitor_bfm APB_MONITOR(APB.monitor_mp);
//apb_agent_bfm APB_AGENT(.APB(APB));
//end

// tbx vif_binding_block
initial begin
  import uvm_pkg::uvm_config_db;
  uvm_config_db #(virtual apb_driver_bfm) C1;
  uvm_config_db #(virtual apb_monitor_bfm) C2;
  C1.set(null, "uvm_test_top", $psprintf("%m.APB_DRIVER") , APB_DRIVER); //APB_AGENT.driver);
  C2.set(null, "uvm_test_top", $psprintf("%m.APB_MONITOR") , APB_MONITOR); // APB_AGENT.monitor);
end

//if(HAS_SPI_AGENT) begin: has_spi_agent
spi_driver_bfm  SPI_DRIVER(SPI.driver_mp);
spi_monitor_bfm SPI_MONITOR(SPI.monitor_mp);
//spi_agent_bfm SPI_AGENT(.SPI(SPI));
//end

// tbx vif_binding_block
initial begin
  import uvm_pkg::uvm_config_db;
  uvm_config_db #(virtual spi_driver_bfm) C1;
  uvm_config_db #(virtual spi_monitor_bfm) C2;
  C1.set(null, "uvm_test_top", $psprintf("%m.SPI_DRIVER") , SPI_DRIVER); //SPI_AGENT.driver);
  C2.set(null, "uvm_test_top", $psprintf("%m.SPI_MONITOR") , SPI_MONITOR); // SPI_AGENT.monitor);
end

// DUT
spi_top DUT(
    // APB Interface:
    .PCLK(PCLK),
    .PRESETN(PRESETn),
    .PSEL(APB.PSEL[0]),
    .PADDR(APB.PADDR[4:0]),
    .PWDATA(APB.PWDATA),
    .PRDATA(APB.PRDATA),
    .PENABLE(APB.PENABLE),
    .PREADY(APB.PREADY),
    .PSLVERR(),
    .PWRITE(APB.PWRITE),
    // Interrupt output
    .IRQ(INTR.IRQ),
    // SPI signals
    .ss_pad_o(SPI.cs),
    .sclk_pad_o(SPI.clk),
    .mosi_pad_o(SPI.mosi),
    .miso_pad_i(SPI.miso)
);


//
// Clock and reset initial blocks:
//
// tbx clkgen
initial begin
  PCLK = 0;
  forever begin
    #10ns PCLK = ~PCLK;
  end
end

// tbx clkgen
initial begin
  PRESETn = 0;
  #80 PRESETn = 1;
end

endmodule: top_hdl
