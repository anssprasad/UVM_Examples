//------------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

module binder();

bind pss
apb_prober probe   (.PCLK(PCLK),
                    .PRESETn(PRESETn),
                    .PADDR(PADDR),
                    .SPI_PRDATA(SPI_PRDATA),
                    .GPIO_PRDATA(GPIO_PRDATA),
                    .ICPIT_PRDATA(ICPIT_PRDATA),
                    .UART_PRDATA(UART_PRDATA),
                    .SPI_PREADY(SPI_PREADY),
                    .GPIO_PREADY(GPIO_PREADY),
                    .ICPIT_PREADY(ICPIT_PREADY),
                    .UART_PREADY(UART_PREADY),
                    .PWDATA(PWDATA),
                    .PSEL(PSEL),
                    .PENABLE(PENABLE),
                    .PWRITE(PWRITE)
                    );

endmodule: binder

