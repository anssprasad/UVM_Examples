//------------------------------------------------------------
//   Copyright 2007-2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//   
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//   
//       http://www.apache.org/licenses/LICENSE-2.0
//   
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

// Package: Simple Bus OVC
// This is the simple_bus OVC.

package simple_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  typedef enum bit { BUS_R, BUS_W } bus_op_t;

  `include "simple_item.svh"
  `include "simple_sequencer.svh"
  `include "simple_driver.svh"
  `include "simple_seq.svh"
  `include "simple_agent.svh"
endpackage
